module 	block_rom(input  [7:0]  addr,
						 output [31:0] data
						 );

parameter ADDR_WIDTH =  8;
parameter DATA_WIDTH =  32;

parameter [0:71][DATA_WIDTH-1:0] ROM = {
			 // empty 'd0
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 // unpressed 'd18
			 32'b00000000000000000000000000000000,
			 32'b00111111111111111111111111111100,
			 32'b01111111111111111111111111111110,
			 32'b01110000000000000000000000001110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01100000000000000000000000000110,
			 32'b01110000000000000000000000001110,
			 32'b01111111111111111111111111111110,
			 32'b00111111111111111111111111111100,
			 32'b00000000000000000000000000000000,
			 // pressed 'd36
			 32'b00001111111111111111111111110000,
			 32'b00111111111111111111111111111100,
			 32'b01111111111111111111111111111110,
			 32'b01111111111111111111111111111110,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b11110000000000000000000000001111,
			 32'b01111111111111111111111111111110,
			 32'b01111111111111111111111111111110,
			 32'b00111111111111111111111111111100,
			 32'b00001111111111111111111111110000,
			 // "notes" 'd54
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00001111111111111111111111110000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000,
			 32'b00000000000000000000000000000000
			 };
			 
assign data = ROM[addr];
endmodule
